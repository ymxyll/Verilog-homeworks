module counter(
    input clk, rst,
    
);


endcase