module beep_beep();




endmodule