module game_top(
    input [15:0]led,

);