module dz_transfer
(
    input clk, cst, dst, rst,//温度高cst0,dst控制点阵显示复位变成蛋,dst=0温度低
    input fail, dz_num,
    output [7:0] row, colg, colr
);

//将dz_num映射为对应的图像输入到dz_show中进行展示
//fail变绿

reg [3:0] num;//传入点阵的控制值
wire [4:0] rand_num;//接收随机数的值

wire [1:0] rand_ans;//决定哪个动物

reg rand_st;//随机数使能

assign rand_ans = rand_num[1:0];//0~3个

//生成随机数，映射到(0,4区间)随机显示动物图像
get_random random
(
    .clk(clk),
    .st(rand_st),
    .rand(rand_num)
);

dz_show dzs
(
    .clk(clk),
    .rst(),
    .fail(fail),
    .st(dst),
    .num(num),
    .row(row),
    .colg(colg),
    .colr(colr)
);//不需要rst

always@(posedge clk or posedge cst or posedge rst)
begin
    if(rst)
    begin
        num <= 4'd0;
    end
    else if(cst)
    begin
        if(dz_num != 5'd16)
        begin
            num <= dz_num / 2;
            rand_st <= 1'd1;
        end
        else
        begin
            rand_st <= 1'd0;
            num <= 4'd8 + rand_ans;
        end            
    end
    else
        num <= num;
end

endmodule