module counter//1s��������2s������
(
    input clk, rst, st,
    output clk_1s, clk_2s
);

endmodule