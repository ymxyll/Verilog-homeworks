//ÿ��ͼ��Ӧһ��״̬�������״̬��Ϣ�Լ��¶���Ϣ(Ҫ����5s��������)����
module eggs_hatch_top
(
    input clk, rst, btn0, sw7, sw0,
    output led0, led2,
    output [7:0] row, colg, colr, seg, dig
);

wire btn0_o;

debounce db
(
    .clk(clk),
    .btn(btn0),
    .btn_o(btn0_o)
);
//��Ҫһ��1scounter������Ҫһ��2scounter


endmodule