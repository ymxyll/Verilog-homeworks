`timescale 1ns/1ns
module get_random_tb();
//input
reg clk, st;