module counter(
    input clk, rst,
    output 
);


endcase