module disp_show(
    input clk, rst, st,
    input 
);