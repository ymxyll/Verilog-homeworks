module counter
(


);

endmodule