//ÿ��ͼ��Ӧһ��״̬�������״̬��Ϣ�Լ��¶���Ϣ(Ҫ����5s��������)����
module eggs_hatch_top(
    input clk, rst, btn0, sw7, sw0,
    output led0, led2,
);