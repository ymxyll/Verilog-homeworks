module counter(
    input clk, rst,
    output reg [7:0] row, colr, colg;
);


endcase