module counter
(
    input clk, rst, st,
    output clk_1s, clk_2s
);

endmodule