module game_top(
    input led[15:0];
    
);