//���Ƶ��
module half_clk(
    input clk,
    output half_clk
);

endmodule