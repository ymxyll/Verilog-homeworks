//���Ƶ��
module half_clk(


);

endmodule