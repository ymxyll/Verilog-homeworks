module counter(
    input clk, rst,
    output wire [7:0] row, colr, colg
);


endmodule