module game_top(
    input clk, start, rst, sure,
    output [15:0]led,//led
    output [7:0] seg,//����
    output [7:0] dig,//λ��
);