module game_top(
    input [15:0]led,//led
    input [7:0] seg,//����
    input [7:0] dig,//λ��
);