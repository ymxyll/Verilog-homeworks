module dz_show(
    input clk,
    input rst,//�߸�λ
    input reg[2:0] num,
    output reg [7:0] row, colr, colg
);

//����״̬��
always @(posedge clk or posedge rst)
begin
    
end

endmodule