`timescale 1ns/1ns
module game_top();
//input