`timescale 1ns/1ns
module dz_counter_tb();
//input
reg clk, rst;
reg [7:0] row, colg, colr;

endmodule