module game_top(
    output [15:0]led,//led
    output [7:0] seg,//����
    output [7:0] dig,//λ��
);