module get_random_tb();
