module dz_show(
    input clk, rst;
    input reg[2:0] num;
    output reg [7:0] row, colr, colg;
);

endmodule