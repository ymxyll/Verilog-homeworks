//ÿ��ͼ��Ӧһ��״̬�������״̬��Ϣ�Լ��¶���Ϣ����
module eggs_hatch_top(
    input clk, rst, btn0, sw7, sw0;
);