module dz_counter_tb();