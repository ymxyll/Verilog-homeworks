module disp_show(
    input clk, rst, st,
    output [7:0] seg, dig
);


endmodule