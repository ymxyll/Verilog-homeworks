`timescale 1ns/1ns
module beep_beep();
//input



endmodule