`timescale 1ns/1ns
module dz_counter_tb();

endmodule