module counter(
    input 
);


endcase